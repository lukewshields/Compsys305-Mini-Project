entity FlappyBird is 
end entity FlappyBird

architecture arc of FlappyBird is
end architecture arc
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

entity pipes1 is 
	port (
	
	);

end entity pipes1

architecture arc of pipes1 is 






end architecture arc